library ieee;
use ieee. std_logic_1164.all;
use ieee. std_logic_arith.all;
use ieee. std_logic_unsigned.all;


package pkg is
	type \1-line-number\ is array (0 to 29) of std_logic_vector(11 downto 0);
	type \26-line-number\ is array(0 to 29) of \1-line-number\;
end package;

package body pkg is
end package body;

library ieee;
use ieee. std_logic_1164.all;
use ieee. std_logic_arith.all;
use ieee. std_logic_unsigned.all;
use ieee. numeric_std.all;

library work;
use work.pkg.all;
 
entity Digit is
	PORT( clk: 		   in std_logic;
			municion:	in integer range 0 to 999;
			digito:		in integer range 0 to 100;
			sprite:		out \26-line-number\
			);
end entity;
 
architecture behavioral of Digit is
	-- Vector 2d space ship sprite
	--type \1-line-ship\ is array (0 to 59) of std_logic_vector(11 downto 0);
	--type \26-line-ship\ is array(0 to 59) of \1-line-ship\;
	signal cero, uno, dos, tres, cuatro, cinco, seis, siete, ocho, nueve, sprite_actual: \26-line-number\;
	signal digSel: integer range 0 to 999;
begin
	cero <= ((x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"));
	uno <= ((x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"));
	dos <= ((x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"));
	tres <= ((x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000"));
	cuatro <= ((x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	cinco <= ((x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"));
	seis <= ((x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"));
	siete <= ((x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	ocho <= ((x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"));
	nueve <= ((x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"000",x"000",x"000",x"000",x"000"));
	
	digSel <= integer((municion/digito) mod 10);
	
	DigitSelection: process(clk, municion)
	begin
		if(clk'event and clk='1')then
			if (digSel = 0) then
				sprite_actual <= cero;
			elsif (digSel = 1) then
				sprite_actual <= uno;
			elsif (digSel = 2) then
				sprite_actual <= dos;
			elsif (digSel = 3) then
				sprite_actual <= tres;
			elsif (digSel = 4) then
				sprite_actual <= cuatro;
			elsif (digSel = 5) then
				sprite_actual <= cinco;
			elsif (digSel = 6) then
				sprite_actual <= seis;
			elsif (digSel = 7) then
				sprite_actual <= siete;
			elsif (digSel = 8) then
				sprite_actual <= ocho;
			elsif (digSel = 9) then
				sprite_actual <= nueve;
			end if;
		end if;
	end process;
	
	sprite <= sprite_actual;

end behavioral;