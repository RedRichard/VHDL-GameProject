library ieee;
use ieee. std_logic_1164.all;
use ieee. std_logic_arith.all;
use ieee. std_logic_unsigned.all;
use ieee.math_real.all;

-- Esta entidad es la encargada de administrar lo que se dibuja de acuerdo a las coordenadas

entity GeneradorVideo is
PORT( control_x:	in integer;
		control_y:	in integer;
		control_fire: in std_logic;
		pos_x:	in integer;
		pos_y:	in integer;
		habilitado:	in std_logic;
		clk:		in std_logic;
		rgb: out std_logic_vector(11 downto 0);
		carril_nave:	in integer range 1 to 7);
end GeneradorVideo;
 
architecture behavioral of GeneradorVideo is
	constant midnight_blue : std_logic_vector(11 downto 0) := x"653";
	constant dark_orchid : std_logic_vector(11 downto 0) := x"225";
	
	constant max_horizontal: integer := 580;
	constant max_vertical: integer := 400;
	
	-- Vector 2d space ship sprite
	type \1-line-ship\ is array (0 to 59) of std_logic_vector(11 downto 0);
	type \26-line-ship\ is array(0 to 59) of \1-line-ship\;
	signal ship, ship_idle1, ship_idle2 : \26-line-ship\;
	
	-- Vector 2d bullet sprite
	type \1-line-bullet\ is array (0 to 3) of std_logic_vector(11 downto 0);
	type \12-line-bullet\ is array (0 to 11) of \1-line-bullet\;
	signal bullet: \12-line-bullet\;
	
	-- Vector 2d meteor sprite
	signal meteor : \26-line-ship\;
	
	-- Contadores reloj
	constant max_count: integer := 25000000;
	constant half_count: integer := 12500000;
	signal count: integer range 0 to max_count;
	
	signal aux_x, aux_y : integer;
	
	-- Reloj sprite
	signal clk_sprite: std_logic := '0';
	
	-- Reloj proyectil
	signal clk_bullet: std_logic := '0';
	
	-- Contador proyectil
	constant max_c_bullet: integer := 10000; -- Esto es lo que controla la velocidad de movimiento del bullet
	signal count_bullet: integer range 0 to max_c_bullet;
	constant max_b_movement: integer := 450;
	signal count_bullet_movement: integer range 0 to max_b_movement;
	signal allow_fire: std_logic := '0';
	
	-- Limites proyectil:
	signal posx_proyectil_izq, posx_proyectil_der, posy_proyectil_superior, posy_proyectil_inferior: integer;
	
	-- Nave:
	signal posx_nave_izq, posx_nave_der, posy_nave_superior, posy_nave_inferior: integer;
	
	-- Corazones:
	type \1-line-heart\ is array (0 to 29) of std_logic_vector(11 downto 0);
	type \30-line-heart\ is array (0 to 29) of \1-line-heart\;
	signal heart: \30-line-heart\;
	
	constant pos_x_cor1 : integer := 585;
	constant pos_x_cor2 : integer := 505;
	constant pos_x_cor3 : integer := 425;
	constant pos_y_cor : integer := 425;
	
	signal aux_x_cor : integer;
	signal aux_y_cor : integer;
	
	signal vida: integer range 0 to 6 := 6;
	
	-- Meteoritos:
	constant posx_met_izq: integer := 10;
	constant posx_met_der: integer := 70;
	constant posy_met_superior: integer := 0;
	constant posy_met_inferior: integer := 60;
	constant spawn_time: integer := 3;
	signal aux_cont_met1: integer range 0 to 3 := 0;
	signal aux_met_x : integer := 0;
	signal aux_met_y : integer := 0;
	
	constant max_m_meteor: integer := 420;		-- posicion mayima en 'y' del meteorito
	constant max_c_meteor: integer := 250000; -- para la velocidad del meteorito (frecuencia)
	signal count_c_meteor: integer := 0;		-- contador de avance en reloj
	signal count_meteor: integer := 0;			-- contador de avance en posicion 'y'
	signal met1_exists: std_logic := '1';		-- indica si existe el meteorito o no
	signal met1_hit: std_logic := '0'; 			-- indica si el meteorito ha golpeado al jugador o no
	
	signal clk_met: std_logic := '0';			-- reloj de velocidad de movimiento. Indica cuando avanzar un pixel.
	
	-- Puntuación
	signal puntuacion: integer range 0 to 999 := 0;
	
begin
	
	ship_idle1 <= ((x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"fff",x"f00",x"f00",x"f00",x"800",x"800",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"555",x"08f",x"555",x"555",x"04b",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"555",x"08f",x"fff",x"fff",x"04b",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"fff",x"fff",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"fff",x"fff",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"aa9",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"aa9",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"aa9",x"aa9",x"555",x"08f",x"08f",x"08f",x"04b",x"332",x"887",x"887",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"887",x"887",x"aa9",x"555",x"fff",x"fff",x"332",x"887",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"f00",x"f00",x"f00",x"800",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"f00",x"f00",x"f00",x"800",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"fff",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"555",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"000",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"555",x"555",x"555",x"555",x"332",x"800",x"800",x"000",x"555",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"000",x"f00",x"f00",x"332",x"332",x"332",x"332",x"332",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"fff",x"555",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"f00",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"fff",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"fff",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"f00",x"555",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"800",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"f00",x"aa9",x"aa9",x"555",x"aa9",x"aa9",x"aa9",x"887",x"800",x"800",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"887",x"887",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"887",x"887",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"aa9",x"aa9",x"887",x"555",x"800",x"800",x"332",x"332",x"555",x"555",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"aa9",x"887",x"887",x"887",x"000",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"000",x"000",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"555",x"aa9",x"887",x"887",x"000",x"ff0",x"000",x"000",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"887",x"800",x"800",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"000",x"880",x"880",x"000",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"555",x"aa9",x"887",x"887",x"000",x"ff0",x"000",x"000",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"887",x"800",x"800",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"000",x"880",x"880",x"000",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"887",x"887",x"555",x"aa9",x"000",x"000",x"ff0",x"000",x"ff0",x"ff0",x"000",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"aa9",x"555",x"800",x"800",x"332",x"555",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"880",x"000",x"000",x"880",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"555",x"555",x"f00",x"aa9",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"887",x"800",x"800",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"555",x"555",x"f00",x"aa9",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"887",x"800",x"800",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"887",x"887",x"887",x"f00",x"f00",x"f00",x"800",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"aa9",x"aa9",x"887",x"555",x"800",x"800",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"800",x"800",x"800",x"800",x"555",x"555",x"332",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"f00",x"f00",x"800",x"800",x"800",x"000",x"000",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"f0f",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"887",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"f0f",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"f00",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"aa9",x"aa9",x"555",x"555",x"555",x"555",x"aa9",x"887",x"887",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"f00",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"aa9",x"aa9",x"555",x"555",x"555",x"555",x"aa9",x"887",x"887",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"332",x"332",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"332",x"332",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	ship_idle2 <= ((x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"fff",x"f00",x"f00",x"f00",x"800",x"800",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"555",x"08f",x"555",x"555",x"04b",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"555",x"08f",x"fff",x"fff",x"04b",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"fff",x"fff",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"fff",x"fff",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"aa9",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"aa9",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"aa9",x"aa9",x"555",x"08f",x"08f",x"08f",x"04b",x"332",x"887",x"887",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"887",x"887",x"aa9",x"555",x"fff",x"fff",x"332",x"887",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"f00",x"f00",x"f00",x"800",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"f00",x"f00",x"f00",x"800",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"fff",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"555",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"000",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"555",x"555",x"555",x"555",x"332",x"800",x"800",x"000",x"555",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"000",x"f00",x"f00",x"332",x"332",x"332",x"332",x"332",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"fff",x"555",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"f00",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"fff",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"fff",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"f00",x"555",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"800",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"f00",x"aa9",x"aa9",x"555",x"aa9",x"aa9",x"aa9",x"887",x"800",x"800",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"887",x"887",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"887",x"887",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"aa9",x"aa9",x"887",x"555",x"800",x"800",x"332",x"332",x"555",x"555",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"aa9",x"887",x"887",x"887",x"000",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"000",x"000",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"555",x"aa9",x"887",x"887",x"000",x"ff0",x"000",x"000",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"887",x"800",x"800",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"000",x"880",x"880",x"000",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"555",x"aa9",x"887",x"887",x"000",x"ff0",x"000",x"000",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"887",x"800",x"800",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"000",x"880",x"880",x"000",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"887",x"887",x"555",x"aa9",x"000",x"000",x"ff0",x"000",x"ff0",x"ff0",x"000",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"aa9",x"555",x"800",x"800",x"332",x"555",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"880",x"000",x"000",x"880",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"555",x"555",x"f00",x"aa9",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"887",x"800",x"800",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"555",x"555",x"f00",x"aa9",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"887",x"800",x"800",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"887",x"887",x"887",x"f00",x"f00",x"f00",x"800",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"aa9",x"aa9",x"887",x"555",x"800",x"800",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"800",x"800",x"800",x"800",x"555",x"555",x"332",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"f00",x"f00",x"800",x"800",x"800",x"000",x"000",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"f0f",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"887",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"f0f",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"f00",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"aa9",x"aa9",x"555",x"555",x"555",x"555",x"aa9",x"887",x"887",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"f00",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"aa9",x"aa9",x"555",x"555",x"555",x"555",x"aa9",x"887",x"887",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"332",x"332",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"332",x"332",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	
	bullet <= ((x"000",x"07f",x"07f",x"000"),(x"07f",x"fff",x"fff",x"07f"),(x"07f",x"fff",x"fff",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"000",x"07f",x"07f",x"000"),(x"000",x"07f",x"07f",x"000"),(x"000",x"07f",x"07f",x"000"));
	
	meteor <= ((x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"000",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"887",x"887",x"887",x"887",x"555",x"332",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"887",x"555",x"555",x"887",x"887",x"aa9",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000"),(x"000",x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000"),(x"000",x"000",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"000",x"000"),(x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"000"),(x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"000"),(x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"000"),(x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"000"),(x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"887",x"887",x"555",x"555",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000"),(x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"000"),(x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"887",x"555",x"555",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000"),(x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"aa9",x"aa9",x"887",x"aa9",x"aa9",x"887",x"555",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332"),(x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"aa9",x"887",x"555",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332"),(x"000",x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"aa9",x"887",x"555",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332"),(x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000"),(x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000"),(x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000"),(x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"000",x"000",x"000"),(x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"332",x"555",x"887",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"aa9",x"aa9",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"332",x"555",x"887",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"887",x"555",x"332",x"555",x"555",x"555",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"555",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"555",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"332",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"887",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"332",x"332",x"332",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"aa9",x"887",x"887",x"887",x"332",x"332",x"555",x"555",x"332",x"332",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"332",x"332",x"332",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	
	heart <= ((x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"fee",x"fee",x"fee",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"fee",x"fee",x"fee",x"fee",x"f00",x"f00",x"f00",x"000"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"fee",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"fee",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"fee",x"fee",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"fee",x"fee",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	
	-- Reloj meteorito:
	ClkMeteor: process(clk)
	begin
		if(clk'event and clk='1')then
			if(count_c_meteor < max_c_meteor)then
				count_c_meteor <= count_c_meteor + 1;
			else
				clk_met <= not clk_met;
				count_c_meteor <= 0;
			end if;
		end if;
	end process;
	
	-- Contador para movimiento de meteorito:
	MeteorMovement: process(clk_met, count_meteor)
	begin
		if(clk_met'event and clk_met = '1')then
			-- if((posy_nave_superior = count_meteor+60) or (posy_nave_superior = count_meteor+30) or (posy_nave_superior = count_meteor) or (posy_nave_inferior = count_meteor + 60) or (posy_nave_inferior = count_meteor + 30) or (posy_nave_inferior = count_meteor)) and (carril_nave = 1) and (met1_exists = '1')then
			if((posy_nave_superior <= count_meteor+60 and posy_nave_superior >= count_meteor) or (posy_nave_inferior <= count_meteor+60 and posy_nave_inferior >= count_meteor))and (carril_nave = 1) and (met1_exists = '1')then	
				vida <= vida - 1; 	-- Aqui quitamos vida cuando se detecta colisión de meteorito
				met1_hit <= '1';
			-- Aquí se destruye el meteorito si choca un proyectil
			elsif (allow_fire = '1') and (posy_proyectil_superior <= posy_met_inferior) and (posx_proyectil_izq >= posx_met_izq and posx_proyectil_der <= posx_met_der) then
				met1_exists <= '0';
				puntuacion <= puntuacion + 1;
			-- Aquí se reinstancia el meteorito después de que se alcanza el límite de la variable count_meteor 
			elsif (met1_exists = '0') and (count_meteor = max_m_meteor) then
				met1_exists <= '1';
				count_meteor <= 0;
			end if;
			if(count_meteor < max_m_meteor) and ((met1_hit = '0') or (met1_exists = '0')) then
				count_meteor <= count_meteor + 1;
			else
				count_meteor <= 0;
				met1_hit <= '0';
			end if;
		end if;
	end process;
	
	-- Reloj para controlar la velocidad de actualización de sprites:
	ClkSpriteUpdateSpeed: process(clk, clk_sprite, count)
	begin
		if(clk'event and clk = '1') then
			if(count = half_count)then
				ship <= ship_idle1;
			end if;
			if(count < max_count)then
				count <= count + 1;
			else
				clk_sprite <= not clk_sprite;
				ship <= ship_idle2;
				count <= 0;
			end if;
		end if;
	end process;
	
	-- Reloj para proyectiles:
	ClkBulletSpeed: process(clk, count_bullet)
	begin
		if(clk'event and clk = '1') then
			if(count_bullet < max_c_bullet)then
				count_bullet <= count_bullet + 1;
			else
				clk_bullet <= not clk_bullet;
				count_bullet <= 0;
			end if;
		end if;
	end process;
	
	-- Contador para movimiento de proyectiles:
	BulletMovement: process(clk_bullet)
	begin
		if(clk_bullet'event and clk_bullet = '1') then
			if(control_fire = '1' and allow_fire = '0')then
				allow_fire <= '1';
				count_bullet_movement <= 0;
			end if;
			if(count_bullet_movement < max_b_movement)then
				count_bullet_movement <= count_bullet_movement + 1;
			else
				allow_fire <= '0';
			end if;
		end if;
	end process;
	
	-- Proceso de dibujo. Test: dibujo de un cuadrado entre 10<=x<=60 y 10<=y<=60
	Draw: process(clk, pos_x, pos_y, habilitado, control_y, control_x)
	begin
		if(clk'event and clk = '1') then
			if(habilitado = '1') then
				-- Cuadrado
				--if((pos_x >= control_x and pos_x <= 60+control_x) and (pos_y >= control_y and pos_y <= 60+control_y))then
				--	rgb <= x"F00";
				
				-- Nave:
				if((pos_x >= control_x+1 and pos_x <= 59+control_x) and (pos_y >= control_y and pos_y <= 60+control_y))then
					aux_x <= pos_x-control_x;
					aux_y <= pos_y-control_y;
					
					rgb <= ship(aux_y)(aux_x);
					
					-- Posiciones de la nave:
					posx_nave_izq <= control_x;
					posx_nave_der <= control_x + 60;
					posy_nave_superior <= control_y;
					posy_nave_inferior <= control_y+60;
					
					-- Esto se utiliza para el disparo del proyectil. Posiciones:
					posx_proyectil_izq <= control_x+28;
					posx_proyectil_der <= 4+control_x+28;
					posy_proyectil_superior <= control_y-count_bullet_movement;
					posy_proyectil_inferior <= 12+control_y-count_bullet_movement;
				-- Proyectil
				elsif ((allow_fire = '1') and (pos_x >= posx_proyectil_izq and pos_x <= posx_proyectil_der) and (pos_y >= posy_proyectil_superior and pos_y <= posy_proyectil_inferior))then
					rgb <= bullet(pos_y)(pos_x);
					
				-- Meteoro 1
				elsif ((met1_exists = '1') and (pos_x >= posx_met_izq and pos_x <= posx_met_der) and (pos_y >= posy_met_superior + count_meteor and pos_y <= posy_met_inferior + count_meteor))then
										
					aux_met_x <= pos_x-posx_met_izq;
					aux_met_y <= pos_y-posy_met_superior-count_meteor;
					rgb <= meteor(aux_met_y)(aux_met_x);
				-- Corazon1
				elsif (vida >= 6) and (pos_x >= pos_x_cor1 and pos_x <= pos_x_cor1+30) and (pos_y >= pos_y_cor and pos_y <= pos_y_cor+30) then
					aux_x_cor <= pos_x - pos_x_cor1;
					aux_y_cor <= pos_y - pos_y_cor;
					rgb <= heart(aux_y_cor)(aux_x_cor);
				-- Corazon2
				elsif (vida >= 4) and (pos_x >= pos_x_cor2 and pos_x <= pos_x_cor2+30) and (pos_y >= pos_y_cor and pos_y <= pos_y_cor+30) then
					aux_x_cor <= pos_x - pos_x_cor2;
					aux_y_cor <= pos_y - pos_y_cor;
					rgb <= heart(aux_y_cor)(aux_x_cor);
				-- Corazon3
				elsif (vida >= 2) and (pos_x >= pos_x_cor3 and pos_x <= pos_x_cor3+30) and (pos_y >= pos_y_cor and pos_y <= pos_y_cor+30) then
					aux_x_cor <= pos_x - pos_x_cor3;
					aux_y_cor <= pos_y - pos_y_cor;
					rgb <= heart(aux_y_cor)(aux_x_cor);
				-- Grid
				elsif (pos_x >= 0 and pos_x <= 2) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= heart(aux_y_cor)(aux_x_cor);
				elsif (pos_x >= 77 and pos_x <= 81) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 157 and pos_x <= 161) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 237 and pos_x <= 241) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 317 and pos_x <= 321) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 397 and pos_x <= 401) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 477 and pos_x <= 481) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 557 and pos_x <= 561) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 637 and pos_x <= 639) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				else
					rgb <= x"000";
				end if;
			else
				rgb <= x"000";
			end if;
		end if;
	end process;
	
	
end behavioral;