library ieee;
use ieee. std_logic_1164.all;
use ieee. std_logic_arith.all;
use ieee. std_logic_unsigned.all;
use ieee.math_real.all;

-- Esta entidad es la encargada de administrar lo que se dibuja de acuerdo a las coordenadas

entity GeneradorVideo is
PORT( control_x:	in integer;
		control_y:	in integer;
		control_fire: in std_logic;
		pos_x:	in integer;
		pos_y:	in integer;
		habilitado:	in std_logic;
		clk:		in std_logic;
		rgb: out std_logic_vector(11 downto 0);
		carril_nave:	in integer range 0 to 8);
end GeneradorVideo;
 
architecture behavioral of GeneradorVideo is
	constant midnight_blue : std_logic_vector(11 downto 0) := x"653";
	constant dark_orchid : std_logic_vector(11 downto 0) := x"225";
	
	constant max_horizontal: integer := 580;
	constant max_vertical: integer := 400;
	
	-- Vector 2d space ship sprite
	type \1-line-ship\ is array (0 to 59) of std_logic_vector(11 downto 0);
	type \26-line-ship\ is array(0 to 59) of \1-line-ship\;
	signal ship, ship_idle1, ship_idle2 : \26-line-ship\;
	
	-- Vector 2d number sprite
	type \1-line-number\ is array (0 to 29) of std_logic_vector(11 downto 0);
	type \26-line-number\ is array(0 to 29) of \1-line-number\;
	signal mun_dig1, mun_dig2: \26-line-number\;
	signal point_dig1, point_dig2, point_dig3: \26-line-number\;
	
	-- Vector 2d bullet sprite
	type \1-line-bullet\ is array (0 to 3) of std_logic_vector(11 downto 0);
	type \12-line-bullet\ is array (0 to 11) of \1-line-bullet\;
	signal bullet: \12-line-bullet\;
	
	-- Vector 2d meteor sprite
	signal meteor : \26-line-ship\;
	
	-- Contadores reloj
	constant max_count: integer := 25000000;
	constant half_count: integer := 12500000;
	signal count: integer range 0 to max_count;
	
	signal aux_x, aux_y : integer;
	
	-- Reloj sprite
	signal clk_sprite: std_logic := '0';
	
	-- Reloj proyectil
	signal clk_bullet: std_logic := '0';
	
	-- Contador proyectil
	constant max_c_bullet: integer := 10000; -- Esto es lo que controla la velocidad de movimiento del bullet
	signal count_bullet: integer range 0 to max_c_bullet;
	constant max_b_movement: integer := 450;
	signal count_bullet_movement: integer range 0 to max_b_movement;
	signal allow_fire: std_logic := '0';
	
	-- Limites proyectil:
	signal posx_proyectil_izq, posx_proyectil_der, posy_proyectil_superior, posy_proyectil_inferior: integer;
	
	-- Nave:
	signal posx_nave_izq, posx_nave_der, posy_nave_superior, posy_nave_inferior: integer;
	
	-- Corazones:
	type \1-line-heart\ is array (0 to 29) of std_logic_vector(11 downto 0);
	type \30-line-heart\ is array (0 to 29) of \1-line-heart\;
	signal heart: \30-line-heart\;
	
	constant pos_x_cor1 : integer := 585;
	constant pos_x_cor2 : integer := 505;
	constant pos_x_cor3 : integer := 425;
	constant pos_y_cor : integer := 425;
	
	signal aux_x_cor : integer;
	signal aux_y_cor : integer;
	
	signal vida: integer range 0 to 999 := 6;
	
	-- Meteoritos:
	--  Meteorito 1:
	constant posx_met1_izq: integer := 10;
	constant posx_met1_der: integer := 70;
	constant posy_met1_superior: integer := -60;
	constant posy_met1_inferior: integer := 0;
	signal aux_met1_x : integer := 0;
	signal aux_met1_y : integer := 0;
	
	signal met1_exists: std_logic;		-- indica si existe el meteorito o no
	signal count_meteor1: integer := 0;			-- contador de avance en posicion 'y'
	signal aux_vida1: integer range 0 to 3; 
	
	--  Meteorito 2:
	constant posx_met2_izq: integer := 90;
	constant posx_met2_der: integer := 150;
	constant posy_met2_superior: integer := -120;
	constant posy_met2_inferior: integer := -60;
	signal aux_met2_x : integer := 0;
	signal aux_met2_y : integer := 0;
	signal aux_vida2: integer range 0 to 3; 
	
	signal met2_exists: std_logic;		-- indica si existe el meteorito o no
	signal count_meteor2: integer := 0;	
	
	--  Meteorito 3:
	constant posx_met3_izq: integer := 170;
	constant posx_met3_der: integer := 230;
	constant posy_met3_superior: integer := -60;
	constant posy_met3_inferior: integer := 0;
	signal aux_met3_x : integer := 0;
	signal aux_met3_y : integer := 0;
	
	signal met3_exists: std_logic;		-- indica si existe el meteorito o no
	signal count_meteor3: integer := 0;			-- contador de avance en posicion 'y'
	signal aux_vida3: integer range 0 to 3; 
	
	--  Meteorito 4:
	constant posx_met4_izq: integer := 250;
	constant posx_met4_der: integer := 310;
	constant posy_met4_superior: integer := -120;
	constant posy_met4_inferior: integer := -60;
	signal aux_met4_x : integer := 0;
	signal aux_met4_y : integer := 0;
	signal aux_vida4: integer range 0 to 3; 
	
	signal met4_exists: std_logic;		-- indica si existe el meteorito o no
	signal count_meteor4: integer := 0;	
	
	--  Meteorito 5:
	constant posx_met5_izq: integer := 330;
	constant posx_met5_der: integer := 390;
	constant posy_met5_superior: integer := -60;
	constant posy_met5_inferior: integer := 0;
	signal aux_met5_x : integer := 0;
	signal aux_met5_y : integer := 0;
	
	signal met5_exists: std_logic;		-- indica si existe el meteorito o no
	signal count_meteor5: integer := 0;			-- contador de avance en posicion 'y'
	signal aux_vida5: integer range 0 to 3;
	
	--  Meteorito 6:
	constant posx_met6_izq: integer := 410;
	constant posx_met6_der: integer := 470;
	constant posy_met6_superior: integer := -120;
	constant posy_met6_inferior: integer := -60;
	signal aux_met6_x : integer := 0;
	signal aux_met6_y : integer := 0;
	signal aux_vida6: integer range 0 to 3; 
	
	signal met6_exists: std_logic;		-- indica si existe el meteorito o no
	signal count_meteor6: integer := 0;	
	
	--  Meteorito 7:
	constant posx_met7_izq: integer := 490;
	constant posx_met7_der: integer := 550;
	constant posy_met7_superior: integer := -60;
	constant posy_met7_inferior: integer := 0;
	signal aux_met7_x : integer := 0;
	signal aux_met7_y : integer := 0;
	
	signal met7_exists: std_logic;		-- indica si existe el meteorito o no
	signal count_meteor7: integer := 0;			-- contador de avance en posicion 'y'
	signal aux_vida7: integer range 0 to 3;
	
	--  Meteorito 8:
	constant posx_met8_izq: integer := 570;
	constant posx_met8_der: integer := 630;
	constant posy_met8_superior: integer := -120;
	constant posy_met8_inferior: integer := -60;
	signal aux_met8_x : integer := 0;
	signal aux_met8_y : integer := 0;
	signal aux_vida8: integer range 0 to 3; 
	
	signal met8_exists: std_logic;		-- indica si existe el meteorito o no
	signal count_meteor8: integer := 0;	
	
	constant max_c_meteor: integer := 250000; -- para la velocidad del meteorito (frecuencia)	
	--constant max_m_meteor: integer := 420;		-- posicion mayima en 'y' del meteorito
	
	--signal count_c_meteor: integer := 0;		-- contador de avance en reloj
	
	
	--signal met1_hit: std_logic := '0'; 			-- indica si el meteorito ha golpeado al jugador o no
	
	--signal clk_met: std_logic := '0';			-- reloj de velocidad de movimiento. Indica cuando avanzar un pixel.
	
	Component Meteorito is
	port(
		new_game: in std_logic;
		num_pantalla: in integer range 0 to 3;
		vida_actual:	in integer range 0 to 3;
		clk: 		in std_logic;
		num_met:		in integer;
		max_c_meteor:	in integer;
		posx_met_der:			in	integer;
		posx_met_izq:			in integer;
		posy_met_inferior:	in integer;
		posy_nave_superior:	in integer;
		posy_nave_inferior:	in integer;
		posy_proyectil_superior:	in integer;
		posx_proyectil_izq:			in integer;
		posx_proyectil_der:			in integer;
		carril_nave:			in integer range 0 to 8;
		allow_fire:				in std_logic;
		aux_vida:				out integer range 0 to 3;
		
		
		met_exists:				out std_logic;
		c_meteor:			out integer
	
	);
	end component;
	
	Component Digit is
	port( clk: 		   in std_logic;
			municion:	in integer range 0 to 999;
			digito:		in integer range 0 to 100;
			sprite:		out \26-line-number\
			);
	end component;
	
	-- Puntuación
	signal puntuacion: integer range 0 to 999 := 000;
	
	-- Munición
	signal municion: integer range 0 to 999 := 10;
	
	signal mun_izq: integer range 0 to 639 := 20;
	--signal mun_der: integer range 0 to 639 := 60;
	--signal mun_arriba: integer range 0 to 479 := 220;
	--signal mun_abajo: integer range 0 to 479 := 260;
	
	--type \1-line-ammo\ is array (0 to 39) of std_logic_vector(11 downto 0);
	--type \40-line-ammo\ is array (0 to 39) of \1-line-ammo\;
	--signal ammo: \40-line-ammo\;
	
	-- Pantalla
	signal num_pantalla: integer range 0 to 3 := 0;
	signal new_game: std_logic;
	--signal clk_aux: std_logic;
	--signal count_aux: integer;
	
	signal add_ammo: std_logic;
	signal allow_add_ammo: std_logic := '0';
	
begin
	new_game <= control_fire;
	
	-- ammo <= ((x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000"),(x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000"),(x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000"),(x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000"),(x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000"),(x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0"),(x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0"),(x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0"),(x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0"),(x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0"),(x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0"),(x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0"),(x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0"),(x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0"),(x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0"),(x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000"),(x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000"),(x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000"),(x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000"),(x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"0f0",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	
	ship_idle1 <= ((x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"fff",x"f00",x"f00",x"f00",x"800",x"800",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"555",x"08f",x"555",x"555",x"04b",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"555",x"08f",x"fff",x"fff",x"04b",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"fff",x"fff",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"fff",x"fff",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"aa9",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"aa9",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"aa9",x"aa9",x"555",x"08f",x"08f",x"08f",x"04b",x"332",x"887",x"887",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"887",x"887",x"aa9",x"555",x"fff",x"fff",x"332",x"887",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"f00",x"f00",x"f00",x"800",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"f00",x"f00",x"f00",x"800",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"fff",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"555",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"000",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"555",x"555",x"555",x"555",x"332",x"800",x"800",x"000",x"555",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"000",x"f00",x"f00",x"332",x"332",x"332",x"332",x"332",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"fff",x"555",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"f00",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"fff",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"fff",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"f00",x"555",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"800",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"f00",x"aa9",x"aa9",x"555",x"aa9",x"aa9",x"aa9",x"887",x"800",x"800",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"887",x"887",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"887",x"887",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"aa9",x"aa9",x"887",x"555",x"800",x"800",x"332",x"332",x"555",x"555",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"aa9",x"887",x"887",x"887",x"000",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"000",x"000",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"555",x"aa9",x"887",x"887",x"000",x"ff0",x"000",x"000",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"887",x"800",x"800",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"000",x"880",x"880",x"000",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"555",x"aa9",x"887",x"887",x"000",x"ff0",x"000",x"000",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"887",x"800",x"800",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"000",x"880",x"880",x"000",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"887",x"887",x"555",x"aa9",x"000",x"000",x"ff0",x"000",x"ff0",x"ff0",x"000",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"aa9",x"555",x"800",x"800",x"332",x"555",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"880",x"000",x"000",x"880",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"555",x"555",x"f00",x"aa9",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"887",x"800",x"800",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"555",x"555",x"f00",x"aa9",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"887",x"800",x"800",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"887",x"887",x"887",x"f00",x"f00",x"f00",x"800",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"aa9",x"aa9",x"887",x"555",x"800",x"800",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"800",x"800",x"800",x"800",x"555",x"555",x"332",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"f00",x"f00",x"800",x"800",x"800",x"000",x"000",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"f0f",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"887",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"f0f",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"f00",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"aa9",x"aa9",x"555",x"555",x"555",x"555",x"aa9",x"887",x"887",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"f00",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"aa9",x"aa9",x"555",x"555",x"555",x"555",x"aa9",x"887",x"887",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"332",x"332",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"332",x"332",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	ship_idle2 <= ((x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"555",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"fff",x"f00",x"f00",x"f00",x"800",x"800",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"555",x"08f",x"555",x"555",x"04b",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"555",x"08f",x"fff",x"fff",x"04b",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"fff",x"fff",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"fff",x"fff",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"887",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"aa9",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"aa9",x"08f",x"08f",x"08f",x"08f",x"04b",x"04b",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"aa9",x"aa9",x"555",x"08f",x"08f",x"08f",x"04b",x"332",x"887",x"887",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"887",x"887",x"aa9",x"555",x"fff",x"fff",x"332",x"887",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"f00",x"f00",x"f00",x"800",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"f00",x"f00",x"f00",x"800",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"fff",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"555",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"000",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"555",x"555",x"555",x"555",x"332",x"800",x"800",x"000",x"555",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"000",x"f00",x"f00",x"332",x"332",x"332",x"332",x"332",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"555",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"fff",x"555",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"f00",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"fff",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"fff",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"555",x"332",x"332",x"f00",x"f00",x"555",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"800",x"800",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"f00",x"f00",x"aa9",x"aa9",x"555",x"aa9",x"aa9",x"aa9",x"887",x"800",x"800",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"887",x"887",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"887",x"887",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"555",x"aa9",x"aa9",x"887",x"555",x"800",x"800",x"332",x"332",x"555",x"555",x"332",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"aa9",x"887",x"887",x"887",x"000",x"887",x"887",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"aa9",x"887",x"800",x"800",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"000",x"000",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"555",x"aa9",x"887",x"887",x"000",x"ff0",x"000",x"000",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"887",x"800",x"800",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"000",x"880",x"880",x"000",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"555",x"aa9",x"887",x"887",x"000",x"ff0",x"000",x"000",x"887",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"887",x"800",x"800",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"000",x"880",x"880",x"000",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"887",x"887",x"555",x"aa9",x"000",x"000",x"ff0",x"000",x"ff0",x"ff0",x"000",x"555",x"555",x"332",x"f00",x"aa9",x"aa9",x"887",x"555",x"555",x"aa9",x"555",x"800",x"800",x"332",x"555",x"332",x"332",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"880",x"000",x"000",x"880",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"555",x"555",x"f00",x"aa9",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"887",x"800",x"800",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"aa9",x"aa9",x"887",x"555",x"555",x"f00",x"aa9",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"887",x"800",x"800",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"887",x"887",x"887",x"f00",x"f00",x"f00",x"800",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"800",x"aa9",x"aa9",x"887",x"aa9",x"aa9",x"887",x"555",x"800",x"800",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"800",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"800",x"800",x"800",x"800",x"555",x"555",x"332",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"f00",x"f00",x"800",x"800",x"800",x"000",x"000",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"f0f",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"887",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"f0f",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"f00",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"aa9",x"aa9",x"555",x"555",x"555",x"555",x"aa9",x"887",x"887",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"f00",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"000",x"aa9",x"aa9",x"555",x"555",x"555",x"555",x"aa9",x"887",x"887",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"f00",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"800",x"800",x"800",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"fff",x"fff",x"f00",x"f00",x"f00",x"f00",x"f00",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"800",x"800",x"800",x"800",x"800",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aa9",x"887",x"887",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"332",x"332",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"332",x"332",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"800",x"800",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"0bf",x"0bf",x"0bf",x"fff",x"fff",x"fff",x"0bf",x"0bf",x"0bf",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"0bf",x"0bf",x"0bf",x"0bf",x"0bf",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"07f",x"07f",x"07f",x"07f",x"07f",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	
	bullet <= ((x"000",x"07f",x"07f",x"000"),(x"07f",x"fff",x"fff",x"07f"),(x"07f",x"fff",x"fff",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"07f",x"0bf",x"0bf",x"07f"),(x"000",x"07f",x"07f",x"000"),(x"000",x"07f",x"07f",x"000"),(x"000",x"07f",x"07f",x"000"));
	
	meteor <= ((x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"000",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"887",x"887",x"887",x"887",x"887",x"555",x"332",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"887",x"555",x"555",x"887",x"887",x"aa9",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000"),(x"000",x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000"),(x"000",x"000",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"000",x"000"),(x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"000"),(x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"000"),(x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"000"),(x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"000"),(x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"887",x"887",x"555",x"555",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"000"),(x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"000"),(x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"887",x"555",x"555",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"000"),(x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"aa9",x"aa9",x"887",x"aa9",x"aa9",x"887",x"555",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332"),(x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"aa9",x"887",x"555",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"555",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332"),(x"000",x"000",x"887",x"aa9",x"aa9",x"887",x"887",x"aa9",x"887",x"555",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332"),(x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000"),(x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000"),(x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000"),(x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"000",x"000",x"000"),(x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"332",x"555",x"887",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"aa9",x"aa9",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"887",x"887",x"555",x"332",x"555",x"887",x"555",x"555",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"887",x"555",x"332",x"555",x"555",x"555",x"332",x"332",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"555",x"555",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"332",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"555",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"555",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"332",x"332",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"555",x"332",x"332",x"332",x"332",x"555",x"332",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"555",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"332",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"332",x"555",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"332",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"332",x"555",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"aa9",x"887",x"332",x"332",x"555",x"555",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"332",x"332",x"332",x"555",x"555",x"555",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"aa9",x"887",x"887",x"887",x"332",x"332",x"555",x"555",x"332",x"332",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"332",x"332",x"332",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"aa9",x"aa9",x"887",x"887",x"887",x"887",x"887",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"887",x"887",x"887",x"887",x"887",x"555",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"555",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	
	heart <= ((x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"fee",x"fee",x"fee",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"fee",x"fee",x"fee",x"fee",x"f00",x"f00",x"f00",x"000"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"fee",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"fee",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"fee",x"fee",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"fee",x"fee",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00"),(x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000"),(x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"f00",x"f00",x"f00",x"f00",x"f00",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	
	Met1: Meteorito port map(new_game, num_pantalla, vida, clk, 0,max_c_meteor, posx_met1_der, posx_met1_izq, posy_met1_inferior, posy_nave_superior, posy_nave_inferior, posy_proyectil_superior, posx_proyectil_izq, posx_proyectil_der,carril_nave,allow_fire, aux_vida1, met1_exists, count_meteor1);
	
	Met2: Meteorito port map(new_game, num_pantalla, vida, clk, 1,max_c_meteor, posx_met2_der, posx_met2_izq, posy_met2_inferior, posy_nave_superior, posy_nave_inferior, posy_proyectil_superior, posx_proyectil_izq, posx_proyectil_der,carril_nave,allow_fire, aux_vida2, met2_exists, count_meteor2);

	Met3: Meteorito port map(new_game, num_pantalla, vida, clk, 2,max_c_meteor, posx_met3_der, posx_met3_izq, posy_met3_inferior, posy_nave_superior, posy_nave_inferior, posy_proyectil_superior, posx_proyectil_izq, posx_proyectil_der,carril_nave,allow_fire, aux_vida3, met3_exists, count_meteor3);
	
	Met4: Meteorito port map(new_game, num_pantalla, vida, clk, 3,max_c_meteor, posx_met4_der, posx_met4_izq, posy_met4_inferior, posy_nave_superior, posy_nave_inferior, posy_proyectil_superior, posx_proyectil_izq, posx_proyectil_der,carril_nave,allow_fire, aux_vida4, met4_exists, count_meteor4);

	Met5: Meteorito port map(new_game, num_pantalla, vida, clk, 4,max_c_meteor, posx_met5_der, posx_met5_izq, posy_met5_inferior, posy_nave_superior, posy_nave_inferior, posy_proyectil_superior, posx_proyectil_izq, posx_proyectil_der,carril_nave,allow_fire, aux_vida5, met5_exists, count_meteor5);

	Met6: Meteorito port map(new_game, num_pantalla, vida, clk, 5,max_c_meteor, posx_met6_der, posx_met6_izq, posy_met6_inferior, posy_nave_superior, posy_nave_inferior, posy_proyectil_superior, posx_proyectil_izq, posx_proyectil_der,carril_nave,allow_fire, aux_vida6, met6_exists, count_meteor6);

	Met7: Meteorito port map(new_game, num_pantalla, vida, clk, 6,max_c_meteor, posx_met7_der, posx_met7_izq, posy_met7_inferior, posy_nave_superior, posy_nave_inferior, posy_proyectil_superior, posx_proyectil_izq, posx_proyectil_der,carril_nave,allow_fire, aux_vida7, met7_exists, count_meteor7);

	Met8: Meteorito port map(new_game, num_pantalla, vida, clk, 7,max_c_meteor, posx_met8_der, posx_met8_izq, posy_met8_inferior, posy_nave_superior, posy_nave_inferior, posy_proyectil_superior, posx_proyectil_izq, posx_proyectil_der,carril_nave,allow_fire, aux_vida8, met8_exists, count_meteor8);

	-- Munición:
	MunDig1: Digit port map(clk, municion, 1,  mun_dig1);
	MunDig2: Digit port map(clk, municion, 10,  mun_dig2);
	
	-- Puntuación:
	PointDig1: Digit port map(clk, puntuacion, 1, point_dig1);
	PointDig2: Digit port map(clk, puntuacion, 10, point_dig2);
	PointDig3: Digit port map(clk, puntuacion, 100, point_dig3);
	
	--Points: process (clk, aux_p1, aux_p2, aux_p3, aux_p4, aux_p5, aux_p6, aux_p7, aux_p8)
	--begin
		--if (clk'event and clk = '1') then
			--if ((aux_p1 = '1') or (aux_p2 = '1') or (aux_p3 = '1') or (aux_p4 = '1') or (aux_p5 = '1') or (aux_p6 = '1') or (aux_p7 = '1') or (aux_p8 = '1')) then
				--puntuacion <= puntuacion + 1;
			--end if;
		--end if;
	--end process;
	
	-- Proceso para cambiar pantalla:
	Pantalla: process (clk)
	begin
		if (clk'event and clk = '1') then
			if (num_pantalla = 0 or num_pantalla = 2) and (control_fire = '1')then
				num_pantalla <= 1;
			elsif (vida = 0) then
				num_pantalla <= 2;
			end if;
		end if;
	end process;
	
	
	-- Proceso para quitar vida: (Ya funciona!!!!)
	Life: process (clk)
	begin
		if (clk'event and clk = '1') then
			if(new_game = '1') and (num_pantalla = 2) then
				vida <= 3;
			end if;
			if (aux_vida1 < vida) then
				vida <= aux_vida1;
			elsif (aux_vida2 < vida) then
				vida <= aux_vida2;
			elsif (aux_vida3 < vida) then
				vida <= aux_vida3;
			elsif (aux_vida4 < vida) then
				vida <= aux_vida4;
			elsif (aux_vida5 < vida) then
				vida <= aux_vida5;
			elsif (aux_vida6 < vida) then
				vida <= aux_vida6;
			elsif (aux_vida7 < vida) then
				vida <= aux_vida7;
			elsif (aux_vida8 < vida) then
				vida <= aux_vida8;
			end if;
		end if;
	end process;
	
	-- Reloj para controlar la velocidad de actualización de sprites de nave y munición adicional:
	ClkSpriteUpdateSpeed: process(clk, clk_sprite, count)
	begin
		if(clk'event and clk = '1') then
			if(count = half_count)then
				ship <= ship_idle1;
				if (mun_izq > 800) then
					mun_izq <= 20;
				else
					mun_izq <= mun_izq + 80;
				end if;
			end if;
			if(count < max_count)then
				count <= count + 1;
			else
				clk_sprite <= not clk_sprite;
				ship <= ship_idle2;
				count <= 0;
			end if;
		end if;
	end process;
	
	-- Detección de obtención de munición adicional y control de munición (cantidades):
	--MoreAmmo: process (clk_bullet)
	--begin
		--if(clk_bullet'event and clk_bullet = '1') then
			--if (new_game = '1') and (num_pantalla = 2) then
				--municion <= 10;
			--end if;
			---if(control_fire = '1' and municion > 0)then
				--municion <= municion - 1; 			-- Reducción de munición
			--end if;
			--if (mun_izq > posx_nave_izq) and (mun_izq < posx_nave_der) and (210 > posy_nave_superior) and (210 < posy_nave_inferior) then
				--municion <= municion + 2;
				--add_ammo <= '1';
			--else
				--add_ammo <= '0';
			--end if;
		--end if;
	--end process;
	
	-- Reloj para proyectiles:
	ClkBulletSpeed: process(clk, count_bullet)
	begin
		if(clk'event and clk = '1') then
			if(count_bullet < max_c_bullet)then
				count_bullet <= count_bullet + 1;
			else
				clk_bullet <= not clk_bullet;
				count_bullet <= 0;
			end if;
		end if;
	end process;
	
	-- Contador para movimiento de proyectiles:
	BulletMovement: process(clk_bullet)
	begin
		if(clk_bullet'event and clk_bullet = '1') then
			if(new_game = '1') and (num_pantalla = 2) then
				puntuacion <= 0;
				--municion <= 10;
			end if;
			if ((allow_add_ammo = '0') and (mun_izq > posx_nave_izq) and (mun_izq < posx_nave_der) and (210 > posy_nave_superior) and (210 < posy_nave_inferior))then
				allow_add_ammo <= '1';
			end if;
			if(control_fire = '1' and allow_fire = '0' and municion > 0)then
				municion <= municion - 1; 			-- Reducción de munición
				puntuacion <= puntuacion + 1;
				allow_fire <= '1';
				count_bullet_movement <= 0;
			elsif (allow_add_ammo = '1') then
				municion <= municion + 1;
				allow_add_ammo <= '0';
			end if;
			if(count_bullet_movement < max_b_movement)then
				count_bullet_movement <= count_bullet_movement + 1;
			else
				allow_fire <= '0';
			end if;
		end if;
	end process;
	
	-- Proceso de dibujo. Test: dibujo de un cuadrado entre 10<=x<=60 y 10<=y<=60
	Draw: process(clk, pos_x, pos_y, habilitado, control_y, control_x)
	begin
		if(clk'event and clk = '1') then
			if(habilitado = '1') and (num_pantalla = 1) then
				-- Nave:
				if((pos_x >= control_x+1 and pos_x <= 59+control_x) and (pos_y >= control_y and pos_y <= 60+control_y))then
					aux_x <= pos_x-control_x;
					aux_y <= pos_y-control_y;
					
					rgb <= ship(aux_y)(aux_x);
					
					-- Posiciones de la nave:
					posx_nave_izq <= control_x;
					posx_nave_der <= control_x + 60;
					posy_nave_superior <= control_y;
					posy_nave_inferior <= control_y+60;
					
					-- Esto se utiliza para el disparo del proyectil. Posiciones:
					posx_proyectil_izq <= control_x+28;
					posx_proyectil_der <= 4+control_x+28;
					posy_proyectil_superior <= control_y-count_bullet_movement;
					posy_proyectil_inferior <= 12+control_y-count_bullet_movement;
					
				-- Proyectil
				elsif ((allow_fire = '1') and (pos_x >= posx_proyectil_izq and pos_x <= posx_proyectil_der) and (pos_y >= posy_proyectil_superior and pos_y <= posy_proyectil_inferior))then
					rgb <= bullet(pos_y)(pos_x);
					
				-- Meteorito 1
				elsif ((met1_exists = '1') and (pos_x >= posx_met1_izq and pos_x <= posx_met1_der) and (pos_y >= posy_met1_superior + count_meteor1 and pos_y <= posy_met1_inferior + count_meteor1))then
										
					aux_met1_x <= pos_x-posx_met1_izq;
					aux_met1_y <= pos_y-posy_met1_superior-count_meteor1;
					rgb <= meteor(aux_met1_y)(aux_met1_x);
				-- Meteorito 2
				elsif ((met2_exists = '1') and (pos_x >= posx_met2_izq and pos_x <= posx_met2_der) and (pos_y >= posy_met2_superior + count_meteor2 and pos_y <= posy_met2_inferior + count_meteor2))then					
					aux_met2_x <= pos_x-posx_met2_izq;
					aux_met2_y <= pos_y-posy_met2_superior-count_meteor2;
					rgb <= meteor(aux_met2_y)(aux_met2_x);
				-- Meteorito 3
				elsif ((met3_exists = '1') and (pos_x >= posx_met3_izq and pos_x <= posx_met3_der) and (pos_y >= posy_met3_superior + count_meteor3 and pos_y <= posy_met3_inferior + count_meteor3))then					
					aux_met3_x <= pos_x-posx_met3_izq;
					aux_met3_y <= pos_y-posy_met3_superior-count_meteor3;
					rgb <= meteor(aux_met3_y)(aux_met3_x);
				-- Meteorito 4
				elsif ((met4_exists = '1') and (pos_x >= posx_met4_izq and pos_x <= posx_met4_der) and (pos_y >= posy_met4_superior + count_meteor4 and pos_y <= posy_met4_inferior + count_meteor4))then					
					aux_met4_x <= pos_x-posx_met4_izq;
					aux_met4_y <= pos_y-posy_met4_superior-count_meteor4;
					rgb <= meteor(aux_met4_y)(aux_met4_x);
				-- Meteorito 5
				elsif ((met5_exists = '1') and (pos_x >= posx_met5_izq and pos_x <= posx_met5_der) and (pos_y >= posy_met5_superior + count_meteor5 and pos_y <= posy_met5_inferior + count_meteor5))then					
					aux_met5_x <= pos_x-posx_met5_izq;
					aux_met5_y <= pos_y-posy_met5_superior-count_meteor5;
					rgb <= meteor(aux_met5_y)(aux_met5_x);
				-- Meteorito 6
				elsif ((met6_exists = '1') and (pos_x >= posx_met6_izq and pos_x <= posx_met6_der) and (pos_y >= posy_met6_superior + count_meteor6 and pos_y <= posy_met6_inferior + count_meteor6))then					
					aux_met6_x <= pos_x-posx_met6_izq;
					aux_met6_y <= pos_y-posy_met6_superior-count_meteor6;
					rgb <= meteor(aux_met6_y)(aux_met6_x);
				-- Meteorito 7
				elsif ((met7_exists = '1') and (pos_x >= posx_met7_izq and pos_x <= posx_met7_der) and (pos_y >= posy_met7_superior + count_meteor7 and pos_y <= posy_met7_inferior + count_meteor7))then					
					aux_met7_x <= pos_x-posx_met7_izq;
					aux_met7_y <= pos_y-posy_met7_superior-count_meteor7;
					rgb <= meteor(aux_met7_y)(aux_met7_x);
				-- Meteorito 8
				elsif ((met8_exists = '1') and (pos_x >= posx_met8_izq and pos_x <= posx_met8_der) and (pos_y >= posy_met8_superior + count_meteor8 and pos_y <= posy_met8_inferior + count_meteor8))then					
					aux_met8_x <= pos_x-posx_met8_izq;
					aux_met8_y <= pos_y-posy_met8_superior-count_meteor8;
					rgb <= meteor(aux_met8_y)(aux_met8_x);
				-- Munición adicional:
				elsif (pos_x >= mun_izq and pos_x <= mun_izq +40) and (pos_y >= 170) and (pos_y <= 210) then
					rgb <= x"FFF";
				-- Corazon1
				elsif (vida = 3) and (pos_x >= pos_x_cor1 and pos_x <= pos_x_cor1+30) and (pos_y >= pos_y_cor and pos_y <= pos_y_cor+30) then
					aux_x_cor <= pos_x - pos_x_cor1;
					aux_y_cor <= pos_y - pos_y_cor;
					rgb <= heart(aux_y_cor)(aux_x_cor);
				-- Corazon2
				elsif (vida >= 2) and (pos_x >= pos_x_cor2 and pos_x <= pos_x_cor2+30) and (pos_y >= pos_y_cor and pos_y <= pos_y_cor+30) then
					aux_x_cor <= pos_x - pos_x_cor2;
					aux_y_cor <= pos_y - pos_y_cor;
					rgb <= heart(aux_y_cor)(aux_x_cor);
				-- Corazon3
				elsif (vida >= 1) and (pos_x >= pos_x_cor3 and pos_x <= pos_x_cor3+30) and (pos_y >= pos_y_cor and pos_y <= pos_y_cor+30) then
					aux_x_cor <= pos_x - pos_x_cor3;
					aux_y_cor <= pos_y - pos_y_cor;
					rgb <= heart(aux_y_cor)(aux_x_cor);
				-- DigitoMunicion1
				elsif (pos_x >= 360 and pos_x <= 390) and (pos_y >= 425 and pos_y <= 455) then
					rgb <= mun_dig1(pos_y - 425)(pos_x - 360);
				-- DigitoMunicion2
				elsif (pos_x >= 330 and pos_x <= 360) and (pos_y >= 425 and pos_y <= 455) then
					rgb <= mun_dig2(pos_y - 425)(pos_x - 330);
				-- DigitoPuntuacion1
				elsif (pos_x >= 200 and pos_x <= 230) and (pos_y >= 425 and pos_y <= 455) then
					rgb <= point_dig1(pos_y - 425)(pos_x - 200);
				-- DigitoPuntuacion2
				elsif (pos_x >= 170 and pos_x <= 200) and (pos_y >= 425 and pos_y <= 455) then
					rgb <= point_dig2(pos_y - 425)(pos_x - 170);
				-- DigitoPuntuacion3
				elsif (pos_x >= 140 and pos_x <= 170) and (pos_y >= 425 and pos_y <= 455) then
					rgb <= point_dig3(pos_y - 425)(pos_x - 140);
				-- Grid
				elsif (pos_x >= 0 and pos_x <= 2) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= heart(aux_y_cor)(aux_x_cor);
				elsif (pos_x >= 77 and pos_x <= 81) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 157 and pos_x <= 161) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 237 and pos_x <= 241) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 317 and pos_x <= 321) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 397 and pos_x <= 401) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 477 and pos_x <= 481) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 557 and pos_x <= 561) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 637 and pos_x <= 639) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				else
					rgb <= x"000";
				end if;
			-- Pantalla de inicio:
			elsif (habilitado = '1') and (num_pantalla = 0) then
				rgb <= x"FFF";
			-- Pantalla de fin de juego:
			elsif (habilitado = '1') and (num_pantalla = 2) then
				rgb <= x"FFF";
			else
				rgb <= x"000";
			end if;
		end if;
	end process;
	
	
end behavioral;