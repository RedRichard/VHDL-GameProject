library ieee;
use ieee. std_logic_1164.all;
use ieee. std_logic_arith.all;
use ieee. std_logic_unsigned.all;
use ieee.math_real.all;

-- Esta entidad es la encargada de administrar lo que se dibuja de acuerdo a las coordenadas

entity GeneradorVideo is
PORT( control_x:	in integer;
		control_y:	in integer;
		pos_x:	in integer;
		pos_y:	in integer;
		habilitado:	in std_logic;
		clk:		in std_logic;
		rgb: out std_logic_vector(11 downto 0));
end GeneradorVideo;
 
architecture behavioral of GeneradorVideo is
	constant midnight_blue : std_logic_vector(11 downto 0) := x"653";
	constant dark_orchid : std_logic_vector(11 downto 0) := x"225";
	
	constant max_horizontal: integer := 580;
	constant max_vertical: integer := 400;
	
	type \1-line\ is array (0 to 59) of std_logic_vector(11 downto 0);
	type \26-line\ is array(0 to 51) of \1-line\;
	signal ship : \26-line\;
	
	signal aux_x, aux_y : integer;
	
begin
	
	ship <= ((x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"200",x"200",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"100",x"400",x"400",x"100",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"300",x"500",x"500",x"300",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"200",x"444",x"655",x"555",x"333",x"200",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"444",x"776",x"777",x"777",x"666",x"444",x"666",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"333",x"666",x"888",x"888",x"988",x"888",x"666",x"333",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"444",x"777",x"888",x"999",x"988",x"888",x"777",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"222",x"444",x"777",x"888",x"444",x"555",x"999",x"777",x"555",x"222",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"322",x"555",x"888",x"999",x"887",x"666",x"999",x"888",x"666",x"333",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"444",x"777",x"999",x"444",x"bbb",x"bbb",x"444",x"999",x"777",x"444",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"444",x"888",x"aaa",x"888",x"ccc",x"ccc",x"777",x"999",x"888",x"444",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"887",x"988",x"aaa",x"ccc",x"ccc",x"aa9",x"aaa",x"666",x"444",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"888",x"444",x"bbb",x"ddd",x"ddd",x"bbb",x"444",x"888",x"666",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"400",x"a00",x"900",x"766",x"999",x"666",x"bbb",x"ddd",x"ddd",x"bbb",x"555",x"a99",x"666",x"900",x"a00",x"400",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"800",x"b00",x"933",x"888",x"777",x"999",x"555",x"666",x"aaa",x"aaa",x"666",x"555",x"aa9",x"666",x"888",x"933",x"b00",x"900",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"988",x"cbb",x"ccc",x"ddd",x"777",x"a99",x"555",x"222",x"887",x"887",x"222",x"555",x"aaa",x"666",x"ddd",x"ccc",x"cbb",x"988",x"533",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"aaa",x"ccc",x"ddd",x"ddd",x"666",x"999",x"555",x"111",x"443",x"443",x"111",x"555",x"aaa",x"666",x"ddd",x"ddd",x"ccc",x"aaa",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"999",x"cbb",x"ddd",x"eee",x"777",x"999",x"777",x"222",x"111",x"111",x"222",x"888",x"aaa",x"666",x"eee",x"ddd",x"cbb",x"999",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"666",x"999",x"baa",x"888",x"877",x"998",x"bbb",x"333",x"110",x"110",x"333",x"bbb",x"998",x"877",x"888",x"baa",x"999",x"666",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"333",x"999",x"bbb",x"ccc",x"ddd",x"baa",x"988",x"bbb",x"555",x"000",x"000",x"445",x"bbb",x"888",x"baa",x"ddd",x"ccc",x"bbb",x"999",x"333",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"444",x"666",x"999",x"ccc",x"edd",x"eee",x"ccc",x"998",x"bbb",x"555",x"222",x"122",x"566",x"aaa",x"888",x"ccc",x"eee",x"edd",x"ccc",x"999",x"666",x"444",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"444",x"666",x"777",x"888",x"ccc",x"eee",x"eee",x"ddd",x"888",x"aaa",x"ccb",x"444",x"444",x"bbb",x"aaa",x"888",x"ddd",x"eee",x"eee",x"ccc",x"888",x"777",x"666",x"444",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"444",x"777",x"777",x"888",x"666",x"ccc",x"eee",x"eee",x"ddd",x"777",x"888",x"bbb",x"555",x"666",x"bbb",x"777",x"666",x"ddd",x"eee",x"eee",x"ccc",x"666",x"888",x"777",x"777",x"444",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"555",x"777",x"888",x"888",x"767",x"666",x"ccc",x"ddd",x"eee",x"eee",x"777",x"888",x"aaa",x"ccc",x"ccc",x"bbb",x"988",x"777",x"eee",x"eee",x"ddd",x"ccc",x"666",x"767",x"888",x"888",x"777",x"555",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"222",x"766",x"777",x"888",x"888",x"888",x"888",x"666",x"bbb",x"ddd",x"eee",x"eee",x"aaa",x"666",x"aaa",x"ccc",x"ccc",x"aaa",x"888",x"aaa",x"eee",x"eee",x"ddd",x"bbb",x"666",x"888",x"888",x"888",x"888",x"777",x"766",x"222",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"222",x"666",x"777",x"888",x"888",x"aaa",x"a99",x"999",x"777",x"bbb",x"aaa",x"eee",x"eee",x"ccc",x"666",x"888",x"bbb",x"bbb",x"bba",x"777",x"ccc",x"eee",x"eee",x"aaa",x"bbb",x"777",x"999",x"a99",x"aaa",x"888",x"888",x"777",x"666",x"222",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"444",x"777",x"888",x"888",x"999",x"aaa",x"988",x"aaa",x"999",x"989",x"aaa",x"ddd",x"eee",x"888",x"888",x"777",x"988",x"bbb",x"baa",x"999",x"777",x"888",x"888",x"eee",x"ddd",x"aaa",x"989",x"999",x"aaa",x"988",x"aaa",x"999",x"888",x"888",x"667",x"444",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"444",x"777",x"888",x"999",x"666",x"a99",x"bbb",x"bbb",x"bbb",x"aaa",x"999",x"777",x"ccc",x"ddd",x"fff",x"ddd",x"bbb",x"999",x"aaa",x"aaa",x"888",x"bbb",x"ddd",x"fff",x"ddd",x"ccc",x"777",x"999",x"aaa",x"bbb",x"bbb",x"bbb",x"a99",x"666",x"999",x"888",x"777",x"444",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"444",x"766",x"888",x"999",x"998",x"a99",x"bbb",x"bbb",x"bbb",x"bbb",x"baa",x"aaa",x"888",x"ddd",x"eee",x"fff",x"edd",x"ccc",x"777",x"999",x"999",x"888",x"ccc",x"edd",x"fff",x"eee",x"ccc",x"888",x"aaa",x"baa",x"bbb",x"bbb",x"bbb",x"bbb",x"a99",x"998",x"999",x"888",x"766",x"444",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"666",x"877",x"777",x"aaa",x"aaa",x"baa",x"bbb",x"ccc",x"bbb",x"cbb",x"bbb",x"aaa",x"aaa",x"666",x"dcc",x"eee",x"fff",x"eee",x"ccc",x"777",x"888",x"888",x"776",x"ccc",x"eee",x"fff",x"eee",x"ccc",x"666",x"aaa",x"aaa",x"bbb",x"cbb",x"bbb",x"ccc",x"bbb",x"baa",x"aaa",x"aaa",x"777",x"877",x"666",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"222",x"665",x"888",x"999",x"aaa",x"aaa",x"bbb",x"bbb",x"ccc",x"ccc",x"ccc",x"ccc",x"ccc",x"bbb",x"aaa",x"666",x"ccc",x"eee",x"fff",x"eee",x"ccc",x"baa",x"888",x"888",x"baa",x"ccc",x"eee",x"fff",x"eee",x"ccc",x"666",x"aaa",x"bbb",x"ccc",x"ccc",x"ccc",x"ccc",x"ccc",x"bbb",x"bbb",x"aaa",x"aaa",x"999",x"888",x"655",x"222",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"222",x"888",x"888",x"999",x"aaa",x"999",x"baa",x"cbb",x"888",x"ccc",x"ddc",x"ccc",x"dcc",x"ccc",x"ccc",x"baa",x"776",x"a99",x"dcc",x"fff",x"eee",x"ccb",x"bbb",x"877",x"777",x"bbb",x"ccb",x"eee",x"fff",x"dcc",x"a99",x"776",x"baa",x"ccc",x"ccc",x"dcc",x"ccc",x"ccc",x"ccc",x"888",x"cbb",x"baa",x"999",x"aaa",x"999",x"888",x"888",x"222",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"400",x"700",x"999",x"aaa",x"888",x"ccb",x"bbb",x"ccc",x"ccc",x"ddd",x"ddd",x"ddd",x"ddd",x"ddd",x"ddd",x"ccc",x"bbb",x"777",x"ccc",x"ddd",x"fff",x"fff",x"ddd",x"ccc",x"777",x"777",x"ccc",x"ddd",x"fff",x"fff",x"ddd",x"ccc",x"777",x"bbb",x"ccc",x"ddd",x"ddd",x"ccc",x"ddd",x"ddd",x"ddd",x"ccc",x"ccc",x"bbb",x"ccb",x"888",x"aaa",x"999",x"700",x"400",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"400",x"700",x"800",x"aaa",x"999",x"bbb",x"ccc",x"ddd",x"999",x"ddd",x"ddd",x"ccc",x"ccc",x"ddd",x"baa",x"ddd",x"ccc",x"bbb",x"766",x"ccc",x"edd",x"fff",x"fff",x"eee",x"ccc",x"999",x"999",x"ccc",x"eee",x"fff",x"fff",x"edd",x"ccc",x"766",x"bbb",x"ccc",x"ddd",x"baa",x"ddd",x"ccc",x"ccc",x"ddd",x"ddd",x"999",x"ddd",x"ccc",x"bbb",x"999",x"aaa",x"800",x"700",x"400",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"600",x"700",x"900",x"700",x"a00",x"cbb",x"ccc",x"dcc",x"aaa",x"ddd",x"ddd",x"ddd",x"ccc",x"ddd",x"ddd",x"ddd",x"ddd",x"ddd",x"bbb",x"766",x"877",x"edd",x"fff",x"fff",x"eee",x"dcc",x"aaa",x"aaa",x"dcc",x"eee",x"ddd",x"ddd",x"edd",x"baa",x"766",x"bbb",x"ddd",x"ddd",x"ddd",x"ddd",x"ddd",x"ccc",x"ddd",x"ddd",x"ddd",x"aaa",x"dcc",x"ccc",x"cbb",x"a00",x"700",x"900",x"700",x"600",x"000",x"000",x"000"),(x"000",x"000",x"500",x"600",x"a00",x"900",x"c00",x"ddd",x"ddd",x"ccc",x"cbb",x"ddd",x"eee",x"eee",x"aaa",x"eee",x"eee",x"eee",x"eee",x"eee",x"ddd",x"bbb",x"888",x"baa",x"ccc",x"fff",x"fff",x"eee",x"ccc",x"aaa",x"aaa",x"ccc",x"eee",x"ddd",x"ddd",x"ccc",x"ccc",x"888",x"bbb",x"ddd",x"eee",x"eee",x"eee",x"eee",x"eee",x"aaa",x"eee",x"eee",x"ddd",x"cbb",x"ccc",x"ddd",x"ddd",x"c00",x"900",x"a00",x"600",x"500",x"000",x"000"),(x"322",x"600",x"800",x"900",x"700",x"c77",x"aaa",x"ddd",x"ddd",x"eee",x"eee",x"eee",x"eee",x"cbb",x"ccc",x"999",x"eee",x"eee",x"eee",x"eee",x"ddd",x"ccc",x"888",x"ccc",x"ddd",x"ddd",x"fff",x"eee",x"ccc",x"99a",x"99a",x"ccc",x"eee",x"ddd",x"bbb",x"ddd",x"ccc",x"777",x"ccc",x"ddd",x"eee",x"eee",x"eee",x"eee",x"999",x"ccc",x"cbb",x"eee",x"eee",x"eee",x"eee",x"ddd",x"ddd",x"aaa",x"c77",x"700",x"900",x"800",x"600",x"222"),(x"400",x"800",x"900",x"700",x"a88",x"bbb",x"999",x"aaa",x"eee",x"eee",x"eee",x"eee",x"cbb",x"ccc",x"ddd",x"ddd",x"eee",x"eee",x"eee",x"eee",x"ddd",x"ccc",x"999",x"888",x"bbb",x"ddd",x"ddd",x"777",x"999",x"767",x"767",x"999",x"777",x"ddd",x"ddd",x"bbb",x"888",x"888",x"ccc",x"ddd",x"eee",x"eee",x"eee",x"eee",x"ddd",x"ddd",x"ccc",x"cbb",x"eee",x"eee",x"eee",x"eee",x"aaa",x"aaa",x"bbb",x"a88",x"700",x"900",x"800",x"400"),(x"300",x"900",x"b00",x"800",x"aaa",x"ddd",x"baa",x"ddd",x"ddd",x"eee",x"888",x"ddd",x"ddd",x"ddd",x"eee",x"eee",x"ccc",x"eee",x"eee",x"eee",x"cbb",x"ccc",x"777",x"999",x"888",x"ddd",x"eee",x"a9a",x"aaa",x"989",x"989",x"aaa",x"a9a",x"eee",x"ddd",x"999",x"999",x"777",x"ccc",x"cbb",x"eee",x"eee",x"eee",x"ccc",x"eee",x"eee",x"ddd",x"ddd",x"ddd",x"888",x"eee",x"ddd",x"ddd",x"baa",x"ddd",x"aaa",x"900",x"b00",x"900",x"300"),(x"ddd",x"600",x"700",x"900",x"cbb",x"cbb",x"eee",x"ddd",x"eee",x"ddd",x"ccc",x"ddd",x"eee",x"edd",x"eee",x"eee",x"ddd",x"eee",x"eee",x"eee",x"bbb",x"ccc",x"777",x"999",x"a99",x"aaa",x"eee",x"ccc",x"aaa",x"999",x"999",x"aaa",x"ccc",x"eee",x"aaa",x"a99",x"999",x"777",x"ccc",x"edd",x"eee",x"eee",x"eee",x"ddd",x"eee",x"eee",x"edd",x"eee",x"ddd",x"ccc",x"ddd",x"eee",x"ddd",x"eee",x"cbb",x"cbb",x"900",x"700",x"600",x"ddd"),(x"000",x"322",x"900",x"a00",x"ccc",x"ddd",x"eee",x"eee",x"ddd",x"ded",x"ddd",x"eee",x"eee",x"eee",x"eee",x"eee",x"ede",x"eee",x"eee",x"eee",x"aaa",x"ccc",x"776",x"ccc",x"dcc",x"999",x"eee",x"ddd",x"bbb",x"a99",x"a99",x"bbb",x"ddd",x"eee",x"999",x"dcc",x"ccc",x"776",x"ccc",x"eee",x"eee",x"eee",x"eee",x"ede",x"eee",x"eee",x"eee",x"eee",x"eee",x"ddd",x"ded",x"ddd",x"eee",x"eee",x"ddd",x"ccc",x"a00",x"600",x"322",x"000"),(x"000",x"000",x"700",x"900",x"a00",x"ddd",x"888",x"ddd",x"eee",x"eee",x"eee",x"fee",x"fff",x"eee",x"fff",x"fff",x"fee",x"efe",x"fff",x"eee",x"bbb",x"cbb",x"777",x"d64",x"ccc",x"999",x"eee",x"ddd",x"bbb",x"aaa",x"aaa",x"bbb",x"ddd",x"eee",x"999",x"ccc",x"d64",x"777",x"cbb",x"eee",x"eee",x"fff",x"efe",x"fee",x"fff",x"fff",x"eee",x"fff",x"fee",x"eee",x"eee",x"eee",x"ddd",x"888",x"ddd",x"a00",x"900",x"700",x"000",x"000"),(x"000",x"000",x"333",x"800",x"a00",x"ccc",x"dcc",x"ddd",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"ddd",x"bbb",x"ccc",x"b33",x"ea9",x"ddd",x"a99",x"aaa",x"999",x"776",x"888",x"888",x"776",x"999",x"aaa",x"a99",x"ddd",x"ea9",x"b33",x"ccc",x"eee",x"ddd",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"eee",x"ddd",x"dcc",x"ccc",x"a00",x"800",x"444",x"000",x"000"),(x"000",x"000",x"000",x"500",x"800",x"ccc",x"ddd",x"ddd",x"ddd",x"ddd",x"eed",x"ddd",x"eee",x"ddd",x"eee",x"eee",x"edd",x"eee",x"ddd",x"ddd",x"ddd",x"ccc",x"d31",x"ea9",x"ddd",x"999",x"ccc",x"bbb",x"aaa",x"999",x"999",x"aaa",x"bbb",x"ccc",x"999",x"ddd",x"ea9",x"d31",x"ccc",x"ddd",x"ddd",x"ddd",x"eee",x"edd",x"eee",x"eee",x"ddd",x"eee",x"ddd",x"eed",x"ddd",x"ddd",x"ddd",x"ddd",x"ccc",x"800",x"500",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"900",x"b00",x"ccc",x"666",x"777",x"887",x"887",x"988",x"999",x"aaa",x"aaa",x"bbb",x"bbb",x"bbb",x"ccb",x"ccc",x"ddd",x"bbb",x"c20",x"ea9",x"cbb",x"baa",x"ddd",x"ccc",x"bbb",x"999",x"999",x"bbb",x"ccc",x"ddd",x"baa",x"cbb",x"ea9",x"c20",x"bbb",x"ddd",x"ccc",x"ccb",x"bbb",x"bbb",x"bbb",x"aaa",x"aaa",x"999",x"988",x"887",x"887",x"777",x"666",x"ccc",x"b00",x"900",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"411",x"800",x"aaa",x"555",x"555",x"666",x"766",x"777",x"777",x"888",x"888",x"999",x"aaa",x"aaa",x"aaa",x"aaa",x"cbb",x"aaa",x"c00",x"ea9",x"dcc",x"bbb",x"eee",x"ccc",x"ccc",x"aaa",x"aaa",x"ccc",x"ccc",x"eee",x"bbb",x"dcc",x"ea9",x"c00",x"aaa",x"cbb",x"aaa",x"aaa",x"aaa",x"aaa",x"999",x"888",x"888",x"777",x"777",x"766",x"666",x"555",x"555",x"aaa",x"800",x"411",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"444",x"332",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"443",x"a00",x"e98",x"ddd",x"bbb",x"ddd",x"dcc",x"ccc",x"aaa",x"aaa",x"ccc",x"dcc",x"ddd",x"bbb",x"ddd",x"e98",x"a00",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"333",x"332",x"322",x"776",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"633",x"e86",x"ddd",x"bab",x"ddd",x"dcc",x"ccc",x"aaa",x"aaa",x"ccc",x"dcc",x"ddd",x"bab",x"ddd",x"e86",x"533",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"333",x"d64",x"edd",x"888",x"444",x"333",x"222",x"111",x"111",x"222",x"333",x"444",x"888",x"edd",x"d64",x"666",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"444",x"ddd",x"777",x"443",x"222",x"222",x"444",x"444",x"222",x"222",x"443",x"777",x"ddd",x"444",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"),(x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"333",x"333",x"111",x"111",x"221",x"333",x"fff",x"fff",x"333",x"111",x"111",x"111",x"333",x"333",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000"));
	
	-- Proceso de dibujo. Test: dibujo de un cuadrado entre 10<=x<=60 y 10<=y<=60
	Draw: process(clk, pos_x, pos_y, habilitado, control_y, control_x)
	begin
		if(clk'event and clk = '1') then
			if(habilitado = '1') then
				-- Cuadrado
				--if((pos_x >= control_x and pos_x <= 60+control_x) and (pos_y >= control_y and pos_y <= 60+control_y))then
				--	rgb <= x"F00";
				
				-- Nave:
				if((pos_x >= control_x and pos_x <= 60+control_x) and (pos_y >= control_y and pos_y <= 52+control_y))then
					aux_x <= max_horizontal-pos_x;
					aux_y <= max_vertical-pos_y;
					
					rgb <= ship(pos_y)(pos_x);
				
				-- Grid
				elsif (pos_x >= 0 and pos_x <= 2) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 77 and pos_x <= 81) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 157 and pos_x <= 161) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 237 and pos_x <= 241) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 317 and pos_x <= 321) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 397 and pos_x <= 401) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 477 and pos_x <= 481) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 557 and pos_x <= 561) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				elsif (pos_x >= 637 and pos_x <= 639) and (pos_y >= 0 and pos_y <= 400) then
					rgb <= x"FFF";
				else
					rgb <= x"000";
				end if;
			else
				rgb <= x"000";
			end if;
		end if;
	end process;
	
	
end behavioral;